// `default_nettype none
//
// module displaySelect(
//     input clk,
//     input [7:0] sw,
//     input switch, 
//     output reg [3:0] nibbleMS,
//     output reg [3:0] nibbleLS
//     );

// 	// add dispNum here

//     // change between dec and hex display
//     always @() begin
//         // if in hex mode, pass switches through
//         if () begin

//         end else begin
//             // determine value to display in most significant display
//             // if (sw >= 7'd90) begin
//             //     nibbleMS = 4'd9;
//             // end else if (sw >= 8'd80) begin
//             //     nibbleMS = 4'd8;
//             // end else if (sw >= 8'd70) begin
//             //     nibbleMS = 4'd7;
//             // end
//             // // calculate least significant digit
//             // nibbleLS =  -  * ;
//         end
//     end
// endmodule
